`timescale 1ns / 1ps

/*
module MBIST_diagnostics (
	diag_scan_in, diag_clk, rst_h, hold_l, debugz, diag_scan_out, diag_monitor
	);

	input diag_scan_in;
	input diag_clk;
	input rst_h;
	input hold_l;
	input debugz;
	output diag_scan_out;
	output diag_monitor;


endmodule
*/
