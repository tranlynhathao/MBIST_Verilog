`timescale 1ns / 1ps

/*
module MBIST_TAP_interface (
	algsel_scan_in, algsel_scan_en, algsel_scan_out, algsel_clock
	);

	input algsel_scan_in;
	input algsel_scan_en;
	input algsel_clock;
	output algsel_scan_out;

endmodule
*/
